.TRAN 1ms 20ms
R1 1 2 1027.796943
R2 3 2 2077.156725
R3 2 5 3115.622524
R4 5 0 4111.059088
R5 5 6 3028.790321
R6 9 7 2029.831647
R7 7 8 1004.549566
Vs 1 0 1.0 ac 1.0 sin(0 6.283185307 1.0k)
Ve 0 9 0V
Hd 5 8 Ve 8145.628939
Gb 6 3 (2,5) 0.007002
C1 6 8 0.000001
.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)
.ic v(6)=8.683696 v(8)=0.000000
.END
